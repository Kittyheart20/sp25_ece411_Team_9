always_comb begin
    mon_itf.valid[0] = dut.monitor_valid;
    mon_itf.order[0] = dut.monitor_order;
    mon_itf.inst[0] = dut.monitor_inst;
    mon_itf.rs1_addr[0] = dut.monitor_rs1_addr;
    mon_itf.rs2_addr[0] = dut.monitor_rs2_addr;
    mon_itf.rs1_rdata[0] = dut.monitor_rs1_rdata;
    mon_itf.rs2_rdata[0] = dut.monitor_rs2_rdata;
    mon_itf.rd_addr[0] = dut.monitor_rd_addr;
    mon_itf.rd_wdata[0] = dut.monitor_rd_wdata;
    mon_itf.pc_rdata[0] = dut.monitor_pc_rdata;
    mon_itf.pc_wdata[0] = dut.monitor_pc_wdata;
    mon_itf.mem_addr[0] = dut.monitor_mem_addr;
    mon_itf.mem_rmask[0] = dut.monitor_mem_rmask;
    mon_itf.mem_wmask[0] = dut.monitor_mem_wmask;
    mon_itf.mem_rdata[0] = dut.monitor_mem_rdata;
    mon_itf.mem_wdata[0] = dut.monitor_mem_wdata;
    mon_itf.valid[1] = '0;
    mon_itf.order[1] = '0;
    mon_itf.inst[1] = '0;
    mon_itf.rs1_addr[1] = '0;
    mon_itf.rs2_addr[1] = '0;
    mon_itf.rs1_rdata[1] = '0;
    mon_itf.rs2_rdata[1] = '0;
    mon_itf.rd_addr[1] = '0;
    mon_itf.rd_wdata[1] = '0;
    mon_itf.pc_rdata[1] = '0;
    mon_itf.pc_wdata[1] = '0;
    mon_itf.mem_addr[1] = '0;
    mon_itf.mem_rmask[1] = '0;
    mon_itf.mem_wmask[1] = '0;
    mon_itf.mem_rdata[1] = '0;
    mon_itf.mem_wdata[1] = '0;
    mon_itf.valid[2] = '0;
    mon_itf.order[2] = '0;
    mon_itf.inst[2] = '0;
    mon_itf.rs1_addr[2] = '0;
    mon_itf.rs2_addr[2] = '0;
    mon_itf.rs1_rdata[2] = '0;
    mon_itf.rs2_rdata[2] = '0;
    mon_itf.rd_addr[2] = '0;
    mon_itf.rd_wdata[2] = '0;
    mon_itf.pc_rdata[2] = '0;
    mon_itf.pc_wdata[2] = '0;
    mon_itf.mem_addr[2] = '0;
    mon_itf.mem_rmask[2] = '0;
    mon_itf.mem_wmask[2] = '0;
    mon_itf.mem_rdata[2] = '0;
    mon_itf.mem_wdata[2] = '0;
    mon_itf.valid[3] = '0;
    mon_itf.order[3] = '0;
    mon_itf.inst[3] = '0;
    mon_itf.rs1_addr[3] = '0;
    mon_itf.rs2_addr[3] = '0;
    mon_itf.rs1_rdata[3] = '0;
    mon_itf.rs2_rdata[3] = '0;
    mon_itf.rd_addr[3] = '0;
    mon_itf.rd_wdata[3] = '0;
    mon_itf.pc_rdata[3] = '0;
    mon_itf.pc_wdata[3] = '0;
    mon_itf.mem_addr[3] = '0;
    mon_itf.mem_rmask[3] = '0;
    mon_itf.mem_wmask[3] = '0;
    mon_itf.mem_rdata[3] = '0;
    mon_itf.mem_wdata[3] = '0;
    mon_itf.valid[4] = '0;
    mon_itf.order[4] = '0;
    mon_itf.inst[4] = '0;
    mon_itf.rs1_addr[4] = '0;
    mon_itf.rs2_addr[4] = '0;
    mon_itf.rs1_rdata[4] = '0;
    mon_itf.rs2_rdata[4] = '0;
    mon_itf.rd_addr[4] = '0;
    mon_itf.rd_wdata[4] = '0;
    mon_itf.pc_rdata[4] = '0;
    mon_itf.pc_wdata[4] = '0;
    mon_itf.mem_addr[4] = '0;
    mon_itf.mem_rmask[4] = '0;
    mon_itf.mem_wmask[4] = '0;
    mon_itf.mem_rdata[4] = '0;
    mon_itf.mem_wdata[4] = '0;
    mon_itf.valid[5] = '0;
    mon_itf.order[5] = '0;
    mon_itf.inst[5] = '0;
    mon_itf.rs1_addr[5] = '0;
    mon_itf.rs2_addr[5] = '0;
    mon_itf.rs1_rdata[5] = '0;
    mon_itf.rs2_rdata[5] = '0;
    mon_itf.rd_addr[5] = '0;
    mon_itf.rd_wdata[5] = '0;
    mon_itf.pc_rdata[5] = '0;
    mon_itf.pc_wdata[5] = '0;
    mon_itf.mem_addr[5] = '0;
    mon_itf.mem_rmask[5] = '0;
    mon_itf.mem_wmask[5] = '0;
    mon_itf.mem_rdata[5] = '0;
    mon_itf.mem_wdata[5] = '0;
    mon_itf.valid[6] = '0;
    mon_itf.order[6] = '0;
    mon_itf.inst[6] = '0;
    mon_itf.rs1_addr[6] = '0;
    mon_itf.rs2_addr[6] = '0;
    mon_itf.rs1_rdata[6] = '0;
    mon_itf.rs2_rdata[6] = '0;
    mon_itf.rd_addr[6] = '0;
    mon_itf.rd_wdata[6] = '0;
    mon_itf.pc_rdata[6] = '0;
    mon_itf.pc_wdata[6] = '0;
    mon_itf.mem_addr[6] = '0;
    mon_itf.mem_rmask[6] = '0;
    mon_itf.mem_wmask[6] = '0;
    mon_itf.mem_rdata[6] = '0;
    mon_itf.mem_wdata[6] = '0;
    mon_itf.valid[7] = '0;
    mon_itf.order[7] = '0;
    mon_itf.inst[7] = '0;
    mon_itf.rs1_addr[7] = '0;
    mon_itf.rs2_addr[7] = '0;
    mon_itf.rs1_rdata[7] = '0;
    mon_itf.rs2_rdata[7] = '0;
    mon_itf.rd_addr[7] = '0;
    mon_itf.rd_wdata[7] = '0;
    mon_itf.pc_rdata[7] = '0;
    mon_itf.pc_wdata[7] = '0;
    mon_itf.mem_addr[7] = '0;
    mon_itf.mem_rmask[7] = '0;
    mon_itf.mem_wmask[7] = '0;
    mon_itf.mem_rdata[7] = '0;
    mon_itf.mem_wdata[7] = '0;
end
