// module top_tb;

//     timeunit 1ps;
//     timeprecision 1ps;

//     int clock_half_period_ps;
//     initial begin
//         $value$plusargs("CLOCK_PERIOD_PS_ECE411=%d", clock_half_period_ps);
//         clock_half_period_ps = clock_half_period_ps / 2;
//     end

//     bit clk;
//     always #(clock_half_period_ps) clk = ~clk;
//     bit rst;

//     initial begin
//         $fsdbDumpfile("dump.fsdb");
//         if ($test$plusargs("NO_DUMP_ALL_ECE411")) begin
//             $fsdbDumpvars(0, dut, "+all");
//             $fsdbDumpoff();
//         end else begin
//             $fsdbDumpvars(0, "+all");
//         end
//         rst = 1'b1;
//         repeat (2) @(posedge clk);
//         rst <= 1'b0;
//     end

//     `include "top_tb.svh"

// endmodule
