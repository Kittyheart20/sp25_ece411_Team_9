module deserializer (
    input   logic           clk,
    input   logic           rst,

    
    output  logic[31:0]      bmem_addr,
    output  logic               bmem_read,
    output  logic               bmem_write,
    output  logic[63:0]      bmem_wdata,
    input   logic               bmem_ready,

    input   logic[31:0]      bmem_raddr,
    input   logic[63:0]      bmem_rdata,
    input   logic               bmem_rvalid,

    output   logic[255:0] dfp_rdata,
    output   logic           dfp_resp
);

endmodule